`default_nettype none

module steieio_sfsm_top (
  input [7:0] io_in,
  output [7:0] io_out
);
    
    wire clk = io_in[0];
    wire reset = io_in[1];
    wire din = io_in[2];
    wire [4:0] gpi = io_in[7:3];

    reg cs;
    reg dout;
    reg [5:0] gpo;

    assign io_out[7:0] = {gpo[5:0],dout,cs};

    reg [32:0] shiftr;
    reg [5:0] countr;

    // external clock is 1000Hz, so need 10 bit counter
    reg [9:0] second_counter;
    reg [3:0] digit;

    always @(posedge clk) begin
        // if reset, set counter to 0
        if (reset) begin
            second_counter <= 0;
            digit <= 0;
        end else begin
            // if up to 16e6
            if (second_counter == MAX_COUNT) begin
                // reset
                second_counter <= 0;

                // increment digit
                digit <= digit + 1'b1;

                // only count from 0 to 9
                if (digit == 9)
                    digit <= 0;

            end else
                // increment counter
                second_counter <= second_counter + 1'b1;
        end
    end

endmodule
